--modp_montymul_V2
--Jack Holly

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity modp_montymul_V2 is
end entity;

architecture beh of modp_montymul_V2 is 

begin 
end architecture; 